module driver_v2_wrapper #(
  parameter HOST_ADDR_WIDTH = 21,
  parameter HOST_DATA_WIDTH = 32,
  parameter HP_ADDR_WIDTH = 48,
  parameter HP_DATA_WIDTH = 128,
  parameter MAIN_ADDR_WIDTH = 34,
  parameter MAIN_DATA_WIDTH = 128,
  parameter SUB_ADDR_WIDTH = 34,
  parameter SUB_DATA_WIDTH = 128
) (
  input wire clk,
  input wire rstn,

  input  wire [HOST_ADDR_WIDTH-1:0]   host_awaddr,
  input  wire [HOST_DATA_WIDTH-1:0]   host_wdata,
  input  wire [HOST_DATA_WIDTH/8-1:0] host_wstrb,
  input  wire [HOST_ADDR_WIDTH-1:0]   host_araddr,
  output wire [HOST_DATA_WIDTH-1:0]   host_rdata,
  input  wire       host_awvalid,
  output wire       host_awready,
  input  wire       host_wvalid,
  output wire       host_wready,
  output wire [1:0] host_bresp,
  output wire       host_bvalid,
  input  wire       host_bready,
  input  wire       host_arvalid,
  output wire       host_arready,
  output wire [1:0] host_rresp,
  output wire       host_rvalid,
  input  wire       host_rready,

  input  wire [HP_ADDR_WIDTH-1:0]   hp_awaddr,
  input  wire [HP_DATA_WIDTH-1:0]   hp_wdata,
  input  wire [HP_DATA_WIDTH/8-1:0] hp_wstrb,
  input  wire [HP_ADDR_WIDTH-1:0]   hp_araddr,
  output wire [HP_DATA_WIDTH-1:0]   hp_rdata,
  input  wire [7:0] hp_awlen,
  input  wire [2:0] hp_awsize,
  input  wire [1:0] hp_awburst,
  input  wire       hp_awvalid,
  output wire       hp_awready,
  input  wire       hp_wlast,
  input  wire       hp_wvalid,
  output wire       hp_wready,
  output wire [1:0] hp_bresp,
  output wire       hp_bvalid,
  input  wire       hp_bready,
  input  wire [7:0] hp_arlen,
  input  wire [2:0] hp_arsize,
  input  wire [1:0] hp_arburst,
  input  wire       hp_arvalid,
  output wire       hp_arready,
  output wire [1:0] hp_rresp,
  output wire       hp_rlast,
  output wire       hp_rvalid,
  input  wire       hp_rready,

  output wire [MAIN_ADDR_WIDTH-1:0]   main_awaddr,
  output wire [MAIN_DATA_WIDTH-1:0]   main_wdata,
  output wire [MAIN_DATA_WIDTH/8-1:0] main_wstrb,
  output wire [MAIN_ADDR_WIDTH-1:0]   main_araddr,
  input  wire [MAIN_DATA_WIDTH-1:0]   main_rdata,
  output wire [7:0] main_awlen,
  output wire [2:0] main_awsize,
  output wire [1:0] main_awburst,
  output wire       main_awvalid,
  input  wire       main_awready,
  output wire       main_wlast,
  output wire       main_wvalid,
  input  wire       main_wready,
  input  wire [1:0] main_bresp,
  input  wire       main_bvalid,
  output wire       main_bready,
  output wire [7:0] main_arlen,
  output wire [2:0] main_arsize,
  output wire [1:0] main_arburst,
  output wire       main_arvalid,
  input  wire       main_arready,
  input  wire [1:0] main_rresp,
  input  wire       main_rlast,
  input  wire       main_rvalid,
  output wire       main_rready,

  output wire [SUB_ADDR_WIDTH-1:0]   sub_awaddr,
  output wire [SUB_DATA_WIDTH-1:0]   sub_wdata,
  output wire [SUB_DATA_WIDTH/8-1:0] sub_wstrb,
  output wire [SUB_ADDR_WIDTH-1:0]   sub_araddr,
  input  wire [SUB_DATA_WIDTH-1:0]   sub_rdata,
  output wire [7:0] sub_awlen,
  output wire [2:0] sub_awsize,
  output wire [1:0] sub_awburst,
  output wire       sub_awvalid,
  input  wire       sub_awready,
  output wire       sub_wlast,
  output wire       sub_wvalid,
  input  wire       sub_wready,
  input  wire [1:0] sub_bresp,
  input  wire       sub_bvalid,
  output wire       sub_bready,
  output wire [7:0] sub_arlen,
  output wire [2:0] sub_arsize,
  output wire [1:0] sub_arburst,
  output wire       sub_arvalid,
  input  wire       sub_arready,
  input  wire [1:0] sub_rresp,
  input  wire       sub_rlast,
  input  wire       sub_rvalid,
  output wire       sub_rready
);

driver_v2 #(
  .HOST_ADDR_WIDTH(HOST_ADDR_WIDTH),
  .HOST_DATA_WIDTH(HOST_DATA_WIDTH),
  .HP_ADDR_WIDTH(HP_ADDR_WIDTH),
  .HP_DATA_WIDTH(HP_DATA_WIDTH),
  .MAIN_ADDR_WIDTH(MAIN_ADDR_WIDTH),
  .MAIN_DATA_WIDTH(MAIN_DATA_WIDTH),
  .SUB_ADDR_WIDTH(SUB_ADDR_WIDTH),
  .SUB_DATA_WIDTH(SUB_DATA_WIDTH)
) driver_v2_inst (
  .clk(clk),
  .rstn(rstn),
  .host_awaddr  (host_awaddr),
  .host_wdata   (host_wdata),
  .host_wstrb   (host_wstrb),
  .host_araddr  (host_araddr),
  .host_rdata   (host_rdata),
  .host_awvalid (host_awvalid),
  .host_awready (host_awready),
  .host_wvalid  (host_wvalid),
  .host_wready  (host_wready),
  .host_bresp   (host_bresp),
  .host_bvalid  (host_bvalid),
  .host_bready  (host_bready),
  .host_arvalid (host_arvalid),
  .host_arready (host_arready),
  .host_rresp   (host_rresp),
  .host_rvalid  (host_rvalid),
  .host_rready  (host_rready),
  .hp_awaddr  (hp_awaddr),
  .hp_wdata   (hp_wdata),
  .hp_wstrb   (hp_wstrb),
  .hp_araddr  (hp_araddr),
  .hp_rdata   (hp_rdata),
  .hp_awlen   (hp_awlen),
  .hp_awsize  (hp_awsize),
  .hp_awburst (hp_awburst),
  .hp_awvalid (hp_awvalid),
  .hp_awready (hp_awready),
  .hp_wlast   (hp_wlast),
  .hp_wvalid  (hp_wvalid),
  .hp_wready  (hp_wready),
  .hp_bresp   (hp_bresp),
  .hp_bvalid  (hp_bvalid),
  .hp_bready  (hp_bready),
  .hp_arlen   (hp_arlen),
  .hp_arsize  (hp_arsize),
  .hp_arburst (hp_arburst),
  .hp_arvalid (hp_arvalid),
  .hp_arready (hp_arready),
  .hp_rresp   (hp_rresp),
  .hp_rlast   (hp_rlast),
  .hp_rvalid  (hp_rvalid),
  .hp_rready  (hp_rready),
  .main_awaddr  (main_awaddr),
  .main_wdata   (main_wdata),
  .main_wstrb   (main_wstrb),
  .main_araddr  (main_araddr),
  .main_rdata   (main_rdata),
  .main_awlen   (main_awlen),
  .main_awsize  (main_awsize),
  .main_awburst (main_awburst),
  .main_awvalid (main_awvalid),
  .main_awready (main_awready),
  .main_wlast   (main_wlast),
  .main_wvalid  (main_wvalid),
  .main_wready  (main_wready),
  .main_bresp   (main_bresp),
  .main_bvalid  (main_bvalid),
  .main_bready  (main_bready),
  .main_arlen   (main_arlen),
  .main_arsize  (main_arsize),
  .main_arburst (main_arburst),
  .main_arvalid (main_arvalid),
  .main_arready (main_arready),
  .main_rresp   (main_rresp),
  .main_rlast   (main_rlast),
  .main_rvalid  (main_rvalid),
  .main_rready  (main_rready),
  .sub_awaddr  (sub_awaddr),
  .sub_wdata   (sub_wdata),
  .sub_wstrb   (sub_wstrb),
  .sub_araddr  (sub_araddr),
  .sub_rdata   (sub_rdata),
  .sub_awlen   (sub_awlen),
  .sub_awsize  (sub_awsize),
  .sub_awburst (sub_awburst),
  .sub_awvalid (sub_awvalid),
  .sub_awready (sub_awready),
  .sub_wlast   (sub_wlast),
  .sub_wvalid  (sub_wvalid),
  .sub_wready  (sub_wready),
  .sub_bresp   (sub_bresp),
  .sub_bvalid  (sub_bvalid),
  .sub_bready  (sub_bready),
  .sub_arlen   (sub_arlen),
  .sub_arsize  (sub_arsize),
  .sub_arburst (sub_arburst),
  .sub_arvalid (sub_arvalid),
  .sub_arready (sub_arready),
  .sub_rresp   (sub_rresp),
  .sub_rlast   (sub_rlast),
  .sub_rvalid  (sub_rvalid),
  .sub_rready  (sub_rready)
);

endmodule