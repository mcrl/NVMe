// PCIE TOP module

module TOP #(
  parameter   PCIE_LINK_WIDTH = 1
) (
  input wire  ddr4_clk_p,
  input wire  sys_reset
);

  

endmodule