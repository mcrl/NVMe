module driver_wrapper #(
  parameter HOST_ADDR_WIDTH = 21,
  parameter HOST_DATA_WIDTH = 32,
  parameter HP_ADDR_WIDTH = 48, // 256TB
  parameter HP_DATA_WIDTH = 128,
  parameter WRSQ_ADDR_WIDTH = 34, // 2MB
  parameter WRSQ_DATA_WIDTH = 512, // 64B = 512b
  parameter WRBUF_ADDR_WIDTH = 34, // 2MB
  parameter WRBUF_DATA_WIDTH = 128, // 128b
  parameter WRSQDB_ADDR_WIDTH = 34, // 4GB
  parameter WRSQDB_DATA_WIDTH = 128, // 128b
  parameter WRCQ_ADDR_WIDTH = 34, // 2MB
  parameter WRCQ_DATA_WIDTH = 128, // 16B = 128b
  parameter WRCQDB_ADDR_WIDTH = 34, // 4GB
  parameter WRCQDB_DATA_WIDTH = 128, // 16B = 128b
  parameter RDSQ_ADDR_WIDTH = 34, // 2MB
  parameter RDSQ_DATA_WIDTH = 512, // 64B = 512b
  parameter RDBUF_ADDR_WIDTH = 34, // 2MB
  parameter RDBUF_DATA_WIDTH = 128, // 128b
  parameter RDSQDB_ADDR_WIDTH = 34, // 4GB
  parameter RDSQDB_DATA_WIDTH = 128, // 128b
  parameter RDCQ_ADDR_WIDTH = 34, // 2MB
  parameter RDCQ_DATA_WIDTH = 128, // 16B = 128b
  parameter RDCQDB_ADDR_WIDTH = 34, // 4GB
  parameter RDCQDB_DATA_WIDTH = 128 // 16B = 128b
) (
  input wire clk,
  input wire rstn,

  // AXIL slave
  input  wire [HOST_ADDR_WIDTH-1:0]   host_awaddr,
  input  wire [HOST_DATA_WIDTH-1:0]   host_wdata,
  input  wire [HOST_DATA_WIDTH/8-1:0] host_wstrb,
  input  wire [HOST_ADDR_WIDTH-1:0]   host_araddr,
  output wire [HOST_DATA_WIDTH-1:0]   host_rdata,
  input  wire       host_awvalid,
  output wire       host_awready,
  input  wire       host_wvalid,
  output wire       host_wready,
  output wire [1:0] host_bresp,
  output wire       host_bvalid,
  input  wire       host_bready,
  input  wire       host_arvalid,
  output wire       host_arready,
  output wire [1:0] host_rresp,
  output wire       host_rvalid,
  input  wire       host_rready,

  // 1 AXIB slave : hp
  // 10 AXIB master : wrsq, wrbuf, wrsqdb, wrcq, wrcqdb, rdsq, rdbuf, rdsqdb, rdcq, rdcqdb

  input  wire [HP_ADDR_WIDTH-1:0]   hp_awaddr,
  input  wire [HP_DATA_WIDTH-1:0]   hp_wdata,
  input  wire [HP_DATA_WIDTH/8-1:0] hp_wstrb,
  input  wire [HP_ADDR_WIDTH-1:0]   hp_araddr,
  output wire [HP_DATA_WIDTH-1:0]   hp_rdata,
  input  wire [7:0] hp_awlen,
  input  wire [2:0] hp_awsize,
  input  wire [1:0] hp_awburst,
  input  wire       hp_awvalid,
  output wire       hp_awready,
  input  wire       hp_wlast,
  input  wire       hp_wvalid,
  output wire       hp_wready,
  output wire [1:0] hp_bresp,
  output wire       hp_bvalid,
  input  wire       hp_bready,
  input  wire [7:0] hp_arlen,
  input  wire [2:0] hp_arsize,
  input  wire [1:0] hp_arburst,
  input  wire       hp_arvalid,
  output wire       hp_arready,
  output wire [1:0] hp_rresp,
  output wire       hp_rlast,
  output wire       hp_rvalid,
  input  wire       hp_rready,

  output wire [WRSQ_ADDR_WIDTH-1:0]   wrsq_awaddr,
  output wire [WRSQ_DATA_WIDTH-1:0]   wrsq_wdata,
  output wire [WRSQ_DATA_WIDTH/8-1:0] wrsq_wstrb,
  output wire [WRSQ_ADDR_WIDTH-1:0]   wrsq_araddr,
  input  wire [WRSQ_DATA_WIDTH-1:0]   wrsq_rdata,
  output wire [7:0] wrsq_awlen,
  output wire [2:0] wrsq_awsize,
  output wire [1:0] wrsq_awburst,
  output wire       wrsq_awvalid,
  input  wire       wrsq_awready,
  output wire       wrsq_wlast,
  output wire       wrsq_wvalid,
  input  wire       wrsq_wready,
  input  wire [1:0] wrsq_bresp,
  input  wire       wrsq_bvalid,
  output wire       wrsq_bready,
  output wire [7:0] wrsq_arlen,
  output wire [2:0] wrsq_arsize,
  output wire [1:0] wrsq_arburst,
  output wire       wrsq_arvalid,
  input  wire       wrsq_arready,
  input  wire [1:0] wrsq_rresp,
  input  wire       wrsq_rlast,
  input  wire       wrsq_rvalid,
  output wire       wrsq_rready,

  output wire [WRBUF_ADDR_WIDTH-1:0]   wrbuf_awaddr,
  output wire [WRBUF_DATA_WIDTH-1:0]   wrbuf_wdata,
  output wire [WRBUF_DATA_WIDTH/8-1:0] wrbuf_wstrb,
  output wire [WRBUF_ADDR_WIDTH-1:0]   wrbuf_araddr,
  input  wire [WRBUF_DATA_WIDTH-1:0]   wrbuf_rdata,
  output wire [7:0] wrbuf_awlen,
  output wire [2:0] wrbuf_awsize,
  output wire [1:0] wrbuf_awburst,
  output wire       wrbuf_awvalid,
  input  wire       wrbuf_awready,
  output wire       wrbuf_wlast,
  output wire       wrbuf_wvalid,
  input  wire       wrbuf_wready,
  input  wire [1:0] wrbuf_bresp,
  input  wire       wrbuf_bvalid,
  output wire       wrbuf_bready,
  output wire [7:0] wrbuf_arlen,
  output wire [2:0] wrbuf_arsize,
  output wire [1:0] wrbuf_arburst,
  output wire       wrbuf_arvalid,
  input  wire       wrbuf_arready,
  input  wire [1:0] wrbuf_rresp,
  input  wire       wrbuf_rlast,
  input  wire       wrbuf_rvalid,
  output wire       wrbuf_rready,

  output wire [WRSQDB_ADDR_WIDTH-1:0]   wrsqdb_awaddr,
  output wire [WRSQDB_DATA_WIDTH-1:0]   wrsqdb_wdata,
  output wire [WRSQDB_DATA_WIDTH/8-1:0] wrsqdb_wstrb,
  output wire [WRSQDB_ADDR_WIDTH-1:0]   wrsqdb_araddr,
  input  wire [WRSQDB_DATA_WIDTH-1:0]   wrsqdb_rdata,
  output wire [7:0] wrsqdb_awlen,
  output wire [2:0] wrsqdb_awsize,
  output wire [1:0] wrsqdb_awburst,
  output wire       wrsqdb_awvalid,
  input  wire       wrsqdb_awready,
  output wire       wrsqdb_wlast,
  output wire       wrsqdb_wvalid,
  input  wire       wrsqdb_wready,
  input  wire [1:0] wrsqdb_bresp,
  input  wire       wrsqdb_bvalid,
  output wire       wrsqdb_bready,
  output wire [7:0] wrsqdb_arlen,
  output wire [2:0] wrsqdb_arsize,
  output wire [1:0] wrsqdb_arburst,
  output wire       wrsqdb_arvalid,
  input  wire       wrsqdb_arready,
  input  wire [1:0] wrsqdb_rresp,
  input  wire       wrsqdb_rlast,
  input  wire       wrsqdb_rvalid,
  output wire       wrsqdb_rready,

  output wire [WRCQ_ADDR_WIDTH-1:0]   wrcq_awaddr,
  output wire [WRCQ_DATA_WIDTH-1:0]   wrcq_wdata,
  output wire [WRCQ_DATA_WIDTH/8-1:0] wrcq_wstrb,
  output wire [WRCQ_ADDR_WIDTH-1:0]   wrcq_araddr,
  input  wire [WRCQ_DATA_WIDTH-1:0]   wrcq_rdata,
  output wire [7:0] wrcq_awlen,
  output wire [2:0] wrcq_awsize,
  output wire [1:0] wrcq_awburst,
  output wire       wrcq_awvalid,
  input  wire       wrcq_awready,
  output wire       wrcq_wlast,
  output wire       wrcq_wvalid,
  input  wire       wrcq_wready,
  input  wire [1:0] wrcq_bresp,
  input  wire       wrcq_bvalid,
  output wire       wrcq_bready,
  output wire [7:0] wrcq_arlen,
  output wire [2:0] wrcq_arsize,
  output wire [1:0] wrcq_arburst,
  output wire       wrcq_arvalid,
  input  wire       wrcq_arready,
  input  wire [1:0] wrcq_rresp,
  input  wire       wrcq_rlast,
  input  wire       wrcq_rvalid,
  output wire       wrcq_rready,

  output wire [WRCQDB_ADDR_WIDTH-1:0]   wrcqdb_awaddr,
  output wire [WRCQDB_DATA_WIDTH-1:0]   wrcqdb_wdata,
  output wire [WRCQDB_DATA_WIDTH/8-1:0] wrcqdb_wstrb,
  output wire [WRCQDB_ADDR_WIDTH-1:0]   wrcqdb_araddr,
  input  wire [WRCQDB_DATA_WIDTH-1:0]   wrcqdb_rdata,
  output wire [7:0] wrcqdb_awlen,
  output wire [2:0] wrcqdb_awsize,
  output wire [1:0] wrcqdb_awburst,
  output wire       wrcqdb_awvalid,
  input  wire       wrcqdb_awready,
  output wire       wrcqdb_wlast,
  output wire       wrcqdb_wvalid,
  input  wire       wrcqdb_wready,
  input  wire [1:0] wrcqdb_bresp,
  input  wire       wrcqdb_bvalid,
  output wire       wrcqdb_bready,
  output wire [7:0] wrcqdb_arlen,
  output wire [2:0] wrcqdb_arsize,
  output wire [1:0] wrcqdb_arburst,
  output wire       wrcqdb_arvalid,
  input  wire       wrcqdb_arready,
  input  wire [1:0] wrcqdb_rresp,
  input  wire       wrcqdb_rlast,
  input  wire       wrcqdb_rvalid,
  output wire       wrcqdb_rready,

  output wire [RDSQ_ADDR_WIDTH-1:0]   rdsq_awaddr,
  output wire [RDSQ_DATA_WIDTH-1:0]   rdsq_wdata,
  output wire [RDSQ_DATA_WIDTH/8-1:0] rdsq_wstrb,
  output wire [RDSQ_ADDR_WIDTH-1:0]   rdsq_araddr,
  input  wire [RDSQ_DATA_WIDTH-1:0]   rdsq_rdata,
  output wire [7:0] rdsq_awlen,
  output wire [2:0] rdsq_awsize,
  output wire [1:0] rdsq_awburst,
  output wire       rdsq_awvalid,
  input  wire       rdsq_awready,
  output wire       rdsq_wlast,
  output wire       rdsq_wvalid,
  input  wire       rdsq_wready,
  input  wire [1:0] rdsq_bresp,
  input  wire       rdsq_bvalid,
  output wire       rdsq_bready,
  output wire [7:0] rdsq_arlen,
  output wire [2:0] rdsq_arsize,
  output wire [1:0] rdsq_arburst,
  output wire       rdsq_arvalid,
  input  wire       rdsq_arready,
  input  wire [1:0] rdsq_rresp,
  input  wire       rdsq_rlast,
  input  wire       rdsq_rvalid,
  output wire       rdsq_rready,

  output wire [RDBUF_ADDR_WIDTH-1:0]   rdbuf_awaddr,
  output wire [RDBUF_DATA_WIDTH-1:0]   rdbuf_wdata,
  output wire [RDBUF_DATA_WIDTH/8-1:0] rdbuf_wstrb,
  output wire [RDBUF_ADDR_WIDTH-1:0]   rdbuf_araddr,
  input  wire [RDBUF_DATA_WIDTH-1:0]   rdbuf_rdata,
  output wire [7:0] rdbuf_awlen,
  output wire [2:0] rdbuf_awsize,
  output wire [1:0] rdbuf_awburst,
  output wire       rdbuf_awvalid,
  input  wire       rdbuf_awready,
  output wire       rdbuf_wlast,
  output wire       rdbuf_wvalid,
  input  wire       rdbuf_wready,
  input  wire [1:0] rdbuf_bresp,
  input  wire       rdbuf_bvalid,
  output wire       rdbuf_bready,
  output wire [7:0] rdbuf_arlen,
  output wire [2:0] rdbuf_arsize,
  output wire [1:0] rdbuf_arburst,
  output wire       rdbuf_arvalid,
  input  wire       rdbuf_arready,
  input  wire [1:0] rdbuf_rresp,
  input  wire       rdbuf_rlast,
  input  wire       rdbuf_rvalid,
  output wire       rdbuf_rready,

  output wire [RDSQDB_ADDR_WIDTH-1:0]   rdsqdb_awaddr,
  output wire [RDSQDB_DATA_WIDTH-1:0]   rdsqdb_wdata,
  output wire [RDSQDB_DATA_WIDTH/8-1:0] rdsqdb_wstrb,
  output wire [RDSQDB_ADDR_WIDTH-1:0]   rdsqdb_araddr,
  input  wire [RDSQDB_DATA_WIDTH-1:0]   rdsqdb_rdata,
  output wire [7:0] rdsqdb_awlen,
  output wire [2:0] rdsqdb_awsize,
  output wire [1:0] rdsqdb_awburst,
  output wire       rdsqdb_awvalid,
  input  wire       rdsqdb_awready,
  output wire       rdsqdb_wlast,
  output wire       rdsqdb_wvalid,
  input  wire       rdsqdb_wready,
  input  wire [1:0] rdsqdb_bresp,
  input  wire       rdsqdb_bvalid,
  output wire       rdsqdb_bready,
  output wire [7:0] rdsqdb_arlen,
  output wire [2:0] rdsqdb_arsize,
  output wire [1:0] rdsqdb_arburst,
  output wire       rdsqdb_arvalid,
  input  wire       rdsqdb_arready,
  input  wire [1:0] rdsqdb_rresp,
  input  wire       rdsqdb_rlast,
  input  wire       rdsqdb_rvalid,
  output wire       rdsqdb_rready,

  output wire [RDCQ_ADDR_WIDTH-1:0]   rdcq_awaddr,
  output wire [RDCQ_DATA_WIDTH-1:0]   rdcq_wdata,
  output wire [RDCQ_DATA_WIDTH/8-1:0] rdcq_wstrb,
  output wire [RDCQ_ADDR_WIDTH-1:0]   rdcq_araddr,
  input  wire [RDCQ_DATA_WIDTH-1:0]   rdcq_rdata,
  output wire [7:0] rdcq_awlen,
  output wire [2:0] rdcq_awsize,
  output wire [1:0] rdcq_awburst,
  output wire       rdcq_awvalid,
  input  wire       rdcq_awready,
  output wire       rdcq_wlast,
  output wire       rdcq_wvalid,
  input  wire       rdcq_wready,
  input  wire [1:0] rdcq_bresp,
  input  wire       rdcq_bvalid,
  output wire       rdcq_bready,
  output wire [7:0] rdcq_arlen,
  output wire [2:0] rdcq_arsize,
  output wire [1:0] rdcq_arburst,
  output wire       rdcq_arvalid,
  input  wire       rdcq_arready,
  input  wire [1:0] rdcq_rresp,
  input  wire       rdcq_rlast,
  input  wire       rdcq_rvalid,
  output wire       rdcq_rready,

  output wire [RDCQDB_ADDR_WIDTH-1:0]   rdcqdb_awaddr,
  output wire [RDCQDB_DATA_WIDTH-1:0]   rdcqdb_wdata,
  output wire [RDCQDB_DATA_WIDTH/8-1:0] rdcqdb_wstrb,
  output wire [RDCQDB_ADDR_WIDTH-1:0]   rdcqdb_araddr,
  input  wire [RDCQDB_DATA_WIDTH-1:0]   rdcqdb_rdata,
  output wire [7:0] rdcqdb_awlen,
  output wire [2:0] rdcqdb_awsize,
  output wire [1:0] rdcqdb_awburst,
  output wire       rdcqdb_awvalid,
  input  wire       rdcqdb_awready,
  output wire       rdcqdb_wlast,
  output wire       rdcqdb_wvalid,
  input  wire       rdcqdb_wready,
  input  wire [1:0] rdcqdb_bresp,
  input  wire       rdcqdb_bvalid,
  output wire       rdcqdb_bready,
  output wire [7:0] rdcqdb_arlen,
  output wire [2:0] rdcqdb_arsize,
  output wire [1:0] rdcqdb_arburst,
  output wire       rdcqdb_arvalid,
  input  wire       rdcqdb_arready,
  input  wire [1:0] rdcqdb_rresp,
  input  wire       rdcqdb_rlast,
  input  wire       rdcqdb_rvalid,
  output wire       rdcqdb_rready
);

driver #(
  .HOST_ADDR_WIDTH(HOST_ADDR_WIDTH),
  .HOST_DATA_WIDTH(HOST_DATA_WIDTH),
  .HP_ADDR_WIDTH(HP_ADDR_WIDTH),
  .HP_DATA_WIDTH(HP_DATA_WIDTH),
  .WRSQ_ADDR_WIDTH(WRSQ_ADDR_WIDTH),
  .WRSQ_DATA_WIDTH(WRSQ_DATA_WIDTH),
  .WRBUF_ADDR_WIDTH(WRBUF_ADDR_WIDTH),
  .WRBUF_DATA_WIDTH(WRBUF_DATA_WIDTH),
  .WRSQDB_ADDR_WIDTH(WRSQDB_ADDR_WIDTH),
  .WRSQDB_DATA_WIDTH(WRSQDB_DATA_WIDTH),
  .WRCQ_ADDR_WIDTH(WRCQ_ADDR_WIDTH),
  .WRCQ_DATA_WIDTH(WRCQ_DATA_WIDTH),
  .WRCQDB_ADDR_WIDTH(WRCQDB_ADDR_WIDTH),
  .WRCQDB_DATA_WIDTH(WRCQDB_DATA_WIDTH),
  .RDSQ_ADDR_WIDTH(RDSQ_ADDR_WIDTH),
  .RDSQ_DATA_WIDTH(RDSQ_DATA_WIDTH),
  .RDBUF_ADDR_WIDTH(RDBUF_ADDR_WIDTH),
  .RDBUF_DATA_WIDTH(RDBUF_DATA_WIDTH),
  .RDSQDB_ADDR_WIDTH(RDSQDB_ADDR_WIDTH),
  .RDSQDB_DATA_WIDTH(RDSQDB_DATA_WIDTH),
  .RDCQ_ADDR_WIDTH(RDCQ_ADDR_WIDTH),
  .RDCQ_DATA_WIDTH(RDCQ_DATA_WIDTH),
  .RDCQDB_ADDR_WIDTH(RDCQDB_ADDR_WIDTH),
  .RDCQDB_DATA_WIDTH(RDCQDB_DATA_WIDTH)
) driver_inst (
  .clk(clk),
  .rstn(rstn),
  .host_awaddr  (host_awaddr),
  .host_wdata   (host_wdata),
  .host_wstrb   (host_wstrb),
  .host_araddr  (host_araddr),
  .host_rdata   (host_rdata),
  .host_awvalid (host_awvalid),
  .host_awready (host_awready),
  .host_wvalid  (host_wvalid),
  .host_wready  (host_wready),
  .host_bresp   (host_bresp),
  .host_bvalid  (host_bvalid),
  .host_bready  (host_bready),
  .host_arvalid (host_arvalid),
  .host_arready (host_arready),
  .host_rresp   (host_rresp),
  .host_rvalid  (host_rvalid),
  .host_rready  (host_rready),
  .hp_awaddr  (hp_awaddr),
  .hp_wdata   (hp_wdata),
  .hp_wstrb   (hp_wstrb),
  .hp_araddr  (hp_araddr),
  .hp_rdata   (hp_rdata),
  .hp_awlen   (hp_awlen),
  .hp_awsize  (hp_awsize),
  .hp_awburst (hp_awburst),
  .hp_awvalid (hp_awvalid),
  .hp_awready (hp_awready),
  .hp_wlast   (hp_wlast),
  .hp_wvalid  (hp_wvalid),
  .hp_wready  (hp_wready),
  .hp_bresp   (hp_bresp),
  .hp_bvalid  (hp_bvalid),
  .hp_bready  (hp_bready),
  .hp_arlen   (hp_arlen),
  .hp_arsize  (hp_arsize),
  .hp_arburst (hp_arburst),
  .hp_arvalid (hp_arvalid),
  .hp_arready (hp_arready),
  .hp_rresp   (hp_rresp),
  .hp_rlast   (hp_rlast),
  .hp_rvalid  (hp_rvalid),
  .hp_rready  (hp_rready),
  .wrsq_awaddr  (wrsq_awaddr),
  .wrsq_wdata   (wrsq_wdata),
  .wrsq_wstrb   (wrsq_wstrb),
  .wrsq_araddr  (wrsq_araddr),
  .wrsq_rdata   (wrsq_rdata),
  .wrsq_awlen   (wrsq_awlen),
  .wrsq_awsize  (wrsq_awsize),
  .wrsq_awburst (wrsq_awburst),
  .wrsq_awvalid (wrsq_awvalid),
  .wrsq_awready (wrsq_awready),
  .wrsq_wlast   (wrsq_wlast),
  .wrsq_wvalid  (wrsq_wvalid),
  .wrsq_wready  (wrsq_wready),
  .wrsq_bresp   (wrsq_bresp),
  .wrsq_bvalid  (wrsq_bvalid),
  .wrsq_bready  (wrsq_bready),
  .wrsq_arlen   (wrsq_arlen),
  .wrsq_arsize  (wrsq_arsize),
  .wrsq_arburst (wrsq_arburst),
  .wrsq_arvalid (wrsq_arvalid),
  .wrsq_arready (wrsq_arready),
  .wrsq_rresp   (wrsq_rresp),
  .wrsq_rlast   (wrsq_rlast),
  .wrsq_rvalid  (wrsq_rvalid),
  .wrsq_rready  (wrsq_rready),
  .wrbuf_awaddr  (wrbuf_awaddr),
  .wrbuf_wdata   (wrbuf_wdata),
  .wrbuf_wstrb   (wrbuf_wstrb),
  .wrbuf_araddr  (wrbuf_araddr),
  .wrbuf_rdata   (wrbuf_rdata),
  .wrbuf_awlen   (wrbuf_awlen),
  .wrbuf_awsize  (wrbuf_awsize),
  .wrbuf_awburst (wrbuf_awburst),
  .wrbuf_awvalid (wrbuf_awvalid),
  .wrbuf_awready (wrbuf_awready),
  .wrbuf_wlast   (wrbuf_wlast),
  .wrbuf_wvalid  (wrbuf_wvalid),
  .wrbuf_wready  (wrbuf_wready),
  .wrbuf_bresp   (wrbuf_bresp),
  .wrbuf_bvalid  (wrbuf_bvalid),
  .wrbuf_bready  (wrbuf_bready),
  .wrbuf_arlen   (wrbuf_arlen),
  .wrbuf_arsize  (wrbuf_arsize),
  .wrbuf_arburst (wrbuf_arburst),
  .wrbuf_arvalid (wrbuf_arvalid),
  .wrbuf_arready (wrbuf_arready),
  .wrbuf_rresp   (wrbuf_rresp),
  .wrbuf_rlast   (wrbuf_rlast),
  .wrbuf_rvalid  (wrbuf_rvalid),
  .wrbuf_rready  (wrbuf_rready),
  .wrsqdb_awaddr  (wrsqdb_awaddr),
  .wrsqdb_wdata   (wrsqdb_wdata),
  .wrsqdb_wstrb   (wrsqdb_wstrb),
  .wrsqdb_araddr  (wrsqdb_araddr),
  .wrsqdb_rdata   (wrsqdb_rdata),
  .wrsqdb_awlen   (wrsqdb_awlen),
  .wrsqdb_awsize  (wrsqdb_awsize),
  .wrsqdb_awburst (wrsqdb_awburst),
  .wrsqdb_awvalid (wrsqdb_awvalid),
  .wrsqdb_awready (wrsqdb_awready),
  .wrsqdb_wlast   (wrsqdb_wlast),
  .wrsqdb_wvalid  (wrsqdb_wvalid),
  .wrsqdb_wready  (wrsqdb_wready),
  .wrsqdb_bresp   (wrsqdb_bresp),
  .wrsqdb_bvalid  (wrsqdb_bvalid),
  .wrsqdb_bready  (wrsqdb_bready),
  .wrsqdb_arlen   (wrsqdb_arlen),
  .wrsqdb_arsize  (wrsqdb_arsize),
  .wrsqdb_arburst (wrsqdb_arburst),
  .wrsqdb_arvalid (wrsqdb_arvalid),
  .wrsqdb_arready (wrsqdb_arready),
  .wrsqdb_rresp   (wrsqdb_rresp),
  .wrsqdb_rlast   (wrsqdb_rlast),
  .wrsqdb_rvalid  (wrsqdb_rvalid),
  .wrsqdb_rready  (wrsqdb_rready),
  .wrcq_awaddr  (wrcq_awaddr),
  .wrcq_wdata   (wrcq_wdata),
  .wrcq_wstrb   (wrcq_wstrb),
  .wrcq_araddr  (wrcq_araddr),
  .wrcq_rdata   (wrcq_rdata),
  .wrcq_awlen   (wrcq_awlen),
  .wrcq_awsize  (wrcq_awsize),
  .wrcq_awburst (wrcq_awburst),
  .wrcq_awvalid (wrcq_awvalid),
  .wrcq_awready (wrcq_awready),
  .wrcq_wlast   (wrcq_wlast),
  .wrcq_wvalid  (wrcq_wvalid),
  .wrcq_wready  (wrcq_wready),
  .wrcq_bresp   (wrcq_bresp),
  .wrcq_bvalid  (wrcq_bvalid),
  .wrcq_bready  (wrcq_bready),
  .wrcq_arlen   (wrcq_arlen),
  .wrcq_arsize  (wrcq_arsize),
  .wrcq_arburst (wrcq_arburst),
  .wrcq_arvalid (wrcq_arvalid),
  .wrcq_arready (wrcq_arready),
  .wrcq_rresp   (wrcq_rresp),
  .wrcq_rlast   (wrcq_rlast),
  .wrcq_rvalid  (wrcq_rvalid),
  .wrcq_rready  (wrcq_rready),
  .wrcqdb_awaddr  (wrcqdb_awaddr),
  .wrcqdb_wdata   (wrcqdb_wdata),
  .wrcqdb_wstrb   (wrcqdb_wstrb),
  .wrcqdb_araddr  (wrcqdb_araddr),
  .wrcqdb_rdata   (wrcqdb_rdata),
  .wrcqdb_awlen   (wrcqdb_awlen),
  .wrcqdb_awsize  (wrcqdb_awsize),
  .wrcqdb_awburst (wrcqdb_awburst),
  .wrcqdb_awvalid (wrcqdb_awvalid),
  .wrcqdb_awready (wrcqdb_awready),
  .wrcqdb_wlast   (wrcqdb_wlast),
  .wrcqdb_wvalid  (wrcqdb_wvalid),
  .wrcqdb_wready  (wrcqdb_wready),
  .wrcqdb_bresp   (wrcqdb_bresp),
  .wrcqdb_bvalid  (wrcqdb_bvalid),
  .wrcqdb_bready  (wrcqdb_bready),
  .wrcqdb_arlen   (wrcqdb_arlen),
  .wrcqdb_arsize  (wrcqdb_arsize),
  .wrcqdb_arburst (wrcqdb_arburst),
  .wrcqdb_arvalid (wrcqdb_arvalid),
  .wrcqdb_arready (wrcqdb_arready),
  .wrcqdb_rresp   (wrcqdb_rresp),
  .wrcqdb_rlast   (wrcqdb_rlast),
  .wrcqdb_rvalid  (wrcqdb_rvalid),
  .wrcqdb_rready  (wrcqdb_rready),
  .rdsq_awaddr  (rdsq_awaddr),
  .rdsq_wdata   (rdsq_wdata),
  .rdsq_wstrb   (rdsq_wstrb),
  .rdsq_araddr  (rdsq_araddr),
  .rdsq_rdata   (rdsq_rdata),
  .rdsq_awlen   (rdsq_awlen),
  .rdsq_awsize  (rdsq_awsize),
  .rdsq_awburst (rdsq_awburst),
  .rdsq_awvalid (rdsq_awvalid),
  .rdsq_awready (rdsq_awready),
  .rdsq_wlast   (rdsq_wlast),
  .rdsq_wvalid  (rdsq_wvalid),
  .rdsq_wready  (rdsq_wready),
  .rdsq_bresp   (rdsq_bresp),
  .rdsq_bvalid  (rdsq_bvalid),
  .rdsq_bready  (rdsq_bready),
  .rdsq_arlen   (rdsq_arlen),
  .rdsq_arsize  (rdsq_arsize),
  .rdsq_arburst (rdsq_arburst),
  .rdsq_arvalid (rdsq_arvalid),
  .rdsq_arready (rdsq_arready),
  .rdsq_rresp   (rdsq_rresp),
  .rdsq_rlast   (rdsq_rlast),
  .rdsq_rvalid  (rdsq_rvalid),
  .rdsq_rready  (rdsq_rready),
  .rdbuf_awaddr  (rdbuf_awaddr),
  .rdbuf_wdata   (rdbuf_wdata),
  .rdbuf_wstrb   (rdbuf_wstrb),
  .rdbuf_araddr  (rdbuf_araddr),
  .rdbuf_rdata   (rdbuf_rdata),
  .rdbuf_awlen   (rdbuf_awlen),
  .rdbuf_awsize  (rdbuf_awsize),
  .rdbuf_awburst (rdbuf_awburst),
  .rdbuf_awvalid (rdbuf_awvalid),
  .rdbuf_awready (rdbuf_awready),
  .rdbuf_wlast   (rdbuf_wlast),
  .rdbuf_wvalid  (rdbuf_wvalid),
  .rdbuf_wready  (rdbuf_wready),
  .rdbuf_bresp   (rdbuf_bresp),
  .rdbuf_bvalid  (rdbuf_bvalid),
  .rdbuf_bready  (rdbuf_bready),
  .rdbuf_arlen   (rdbuf_arlen),
  .rdbuf_arsize  (rdbuf_arsize),
  .rdbuf_arburst (rdbuf_arburst),
  .rdbuf_arvalid (rdbuf_arvalid),
  .rdbuf_arready (rdbuf_arready),
  .rdbuf_rresp   (rdbuf_rresp),
  .rdbuf_rlast   (rdbuf_rlast),
  .rdbuf_rvalid  (rdbuf_rvalid),
  .rdbuf_rready  (rdbuf_rready),
  .rdsqdb_awaddr  (rdsqdb_awaddr),
  .rdsqdb_wdata   (rdsqdb_wdata),
  .rdsqdb_wstrb   (rdsqdb_wstrb),
  .rdsqdb_araddr  (rdsqdb_araddr),
  .rdsqdb_rdata   (rdsqdb_rdata),
  .rdsqdb_awlen   (rdsqdb_awlen),
  .rdsqdb_awsize  (rdsqdb_awsize),
  .rdsqdb_awburst (rdsqdb_awburst),
  .rdsqdb_awvalid (rdsqdb_awvalid),
  .rdsqdb_awready (rdsqdb_awready),
  .rdsqdb_wlast   (rdsqdb_wlast),
  .rdsqdb_wvalid  (rdsqdb_wvalid),
  .rdsqdb_wready  (rdsqdb_wready),
  .rdsqdb_bresp   (rdsqdb_bresp),
  .rdsqdb_bvalid  (rdsqdb_bvalid),
  .rdsqdb_bready  (rdsqdb_bready),
  .rdsqdb_arlen   (rdsqdb_arlen),
  .rdsqdb_arsize  (rdsqdb_arsize),
  .rdsqdb_arburst (rdsqdb_arburst),
  .rdsqdb_arvalid (rdsqdb_arvalid),
  .rdsqdb_arready (rdsqdb_arready),
  .rdsqdb_rresp   (rdsqdb_rresp),
  .rdsqdb_rlast   (rdsqdb_rlast),
  .rdsqdb_rvalid  (rdsqdb_rvalid),
  .rdsqdb_rready  (rdsqdb_rready),
  .rdcq_awaddr  (rdcq_awaddr),
  .rdcq_wdata   (rdcq_wdata),
  .rdcq_wstrb   (rdcq_wstrb),
  .rdcq_araddr  (rdcq_araddr),
  .rdcq_rdata   (rdcq_rdata),
  .rdcq_awlen   (rdcq_awlen),
  .rdcq_awsize  (rdcq_awsize),
  .rdcq_awburst (rdcq_awburst),
  .rdcq_awvalid (rdcq_awvalid),
  .rdcq_awready (rdcq_awready),
  .rdcq_wlast   (rdcq_wlast),
  .rdcq_wvalid  (rdcq_wvalid),
  .rdcq_wready  (rdcq_wready),
  .rdcq_bresp   (rdcq_bresp),
  .rdcq_bvalid  (rdcq_bvalid),
  .rdcq_bready  (rdcq_bready),
  .rdcq_arlen   (rdcq_arlen),
  .rdcq_arsize  (rdcq_arsize),
  .rdcq_arburst (rdcq_arburst),
  .rdcq_arvalid (rdcq_arvalid),
  .rdcq_arready (rdcq_arready),
  .rdcq_rresp   (rdcq_rresp),
  .rdcq_rlast   (rdcq_rlast),
  .rdcq_rvalid  (rdcq_rvalid),
  .rdcq_rready  (rdcq_rready),
  .rdcqdb_awaddr  (rdcqdb_awaddr),
  .rdcqdb_wdata   (rdcqdb_wdata),
  .rdcqdb_wstrb   (rdcqdb_wstrb),
  .rdcqdb_araddr  (rdcqdb_araddr),
  .rdcqdb_rdata   (rdcqdb_rdata),
  .rdcqdb_awlen   (rdcqdb_awlen),
  .rdcqdb_awsize  (rdcqdb_awsize),
  .rdcqdb_awburst (rdcqdb_awburst),
  .rdcqdb_awvalid (rdcqdb_awvalid),
  .rdcqdb_awready (rdcqdb_awready),
  .rdcqdb_wlast   (rdcqdb_wlast),
  .rdcqdb_wvalid  (rdcqdb_wvalid),
  .rdcqdb_wready  (rdcqdb_wready),
  .rdcqdb_bresp   (rdcqdb_bresp),
  .rdcqdb_bvalid  (rdcqdb_bvalid),
  .rdcqdb_bready  (rdcqdb_bready),
  .rdcqdb_arlen   (rdcqdb_arlen),
  .rdcqdb_arsize  (rdcqdb_arsize),
  .rdcqdb_arburst (rdcqdb_arburst),
  .rdcqdb_arvalid (rdcqdb_arvalid),
  .rdcqdb_arready (rdcqdb_arready),
  .rdcqdb_rresp   (rdcqdb_rresp),
  .rdcqdb_rlast   (rdcqdb_rlast),
  .rdcqdb_rvalid  (rdcqdb_rvalid),
  .rdcqdb_rready  (rdcqdb_rready)
);

endmodule