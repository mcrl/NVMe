// HP: AXIB slave to kernel
// LP: AXIL slave to kernel
// NL: AXIL master to NVMe
// NM: AXIB master to NVMe
// NS: AXIB slave to NVMe
module driver_wrapper #(
  parameter HP_ADDR_WIDTH = 48,
  parameter HP_DATA_WIDTH = 128,
  parameter LP_ADDR_WIDTH = 32,
  parameter LP_DATA_WIDTH = 32,
  parameter NL_ADDR_WIDTH = 32,
  parameter NL_DATA_WIDTH = 32,
  parameter NM_ADDR_WIDTH = 32,
  parameter NM_DATA_WIDTH = 128,
  parameter NS_ID_WIDTH = 4, // required by DMA IP; otherwise block design emit error
  parameter NS_ADDR_WIDTH = 32,
  parameter NS_DATA_WIDTH = 128,
  parameter SQ_ADDR_WIDTH = 9,
  parameter SQ_DATA_WIDTH = 512
) (
  input wire clk,
  input wire rstn,

  // AXIB slave
  input  wire [HP_ADDR_WIDTH-1:0]   hp_awaddr,
  input  wire [HP_DATA_WIDTH-1:0]   hp_wdata,
  input  wire [HP_DATA_WIDTH/8-1:0] hp_wstrb,
  input  wire [HP_ADDR_WIDTH-1:0]   hp_araddr,
  output wire [HP_DATA_WIDTH-1:0]   hp_rdata,
  input  wire [7:0] hp_awlen,
  input  wire [2:0] hp_awsize,
  input  wire [1:0] hp_awburst,
  input  wire       hp_awvalid,
  output wire       hp_awready,
  input  wire       hp_wlast,
  input  wire       hp_wvalid,
  output wire       hp_wready,
  output wire [1:0] hp_bresp,
  output wire       hp_bvalid,
  input  wire       hp_bready,
  input  wire [7:0] hp_arlen,
  input  wire [2:0] hp_arsize,
  input  wire [1:0] hp_arburst,
  input  wire       hp_arvalid,
  output wire       hp_arready,
  output wire [1:0] hp_rresp,
  output wire       hp_rlast,
  output wire       hp_rvalid,
  input  wire       hp_rready,

  // AXIL slave
  input  wire [LP_ADDR_WIDTH-1:0]   lp_awaddr,
  input  wire [LP_DATA_WIDTH-1:0]   lp_wdata,
  input  wire [LP_DATA_WIDTH/8-1:0] lp_wstrb,
  input  wire [LP_ADDR_WIDTH-1:0]   lp_araddr,
  output wire [LP_DATA_WIDTH-1:0]   lp_rdata,
  input  wire       lp_awvalid,
  output wire       lp_awready,
  input  wire       lp_wvalid,
  output wire       lp_wready,
  output wire [1:0] lp_bresp,
  output wire       lp_bvalid,
  input  wire       lp_bready,
  input  wire       lp_arvalid,
  output wire       lp_arready,
  output wire [1:0] lp_rresp,
  output wire       lp_rvalid,
  input  wire       lp_rready,

  // AXIL master
  output wire [NL_ADDR_WIDTH-1:0]   nl_awaddr,
  output wire [NL_DATA_WIDTH-1:0]   nl_wdata,
  output wire [NL_DATA_WIDTH/8-1:0] nl_wstrb,
  output wire [NL_ADDR_WIDTH-1:0]   nl_araddr,
  input  wire [NL_DATA_WIDTH-1:0]   nl_rdata,
  output wire       nl_awvalid,
  input  wire       nl_awready,
  output wire       nl_wvalid,
  input  wire       nl_wready,
  input  wire [1:0] nl_bresp,
  input  wire       nl_bvalid,
  output wire       nl_bready,
  output wire       nl_arvalid,
  input  wire       nl_arready,
  input  wire [1:0] nl_rresp,
  input  wire       nl_rvalid,
  output wire       nl_rready,

  // AXIB master
  output wire [NM_ADDR_WIDTH-1:0]   nm_awaddr,
  output wire [NM_DATA_WIDTH-1:0]   nm_wdata,
  output wire [NM_DATA_WIDTH/8-1:0] nm_wstrb,
  output wire [NM_ADDR_WIDTH-1:0]   nm_araddr,
  input  wire [NM_DATA_WIDTH-1:0]   nm_rdata,
  output wire [7:0] nm_awlen,
  output wire [2:0] nm_awsize,
  output wire [1:0] nm_awburst,
  output wire       nm_awvalid,
  input  wire       nm_awready,
  output wire       nm_wlast,
  output wire       nm_wvalid,
  input  wire       nm_wready,
  input  wire [1:0] nm_bresp,
  input  wire       nm_bvalid,
  output wire       nm_bready,
  output wire [7:0] nm_arlen,
  output wire [2:0] nm_arsize,
  output wire [1:0] nm_arburst,
  output wire       nm_arvalid,
  input  wire       nm_arready,
  input  wire [1:0] nm_rresp,
  input  wire       nm_rlast,
  input  wire       nm_rvalid,
  output wire       nm_rready,

  // AXIB slave
  input  wire [NS_ID_WIDTH-1:0]     ns_awid,
  input  wire [NS_ADDR_WIDTH-1:0]   ns_awaddr,
  input  wire [NS_DATA_WIDTH-1:0]   ns_wdata,
  input  wire [NS_DATA_WIDTH/8-1:0] ns_wstrb,
  output wire [NS_ID_WIDTH-1:0]     ns_bid,
  input  wire [NS_ID_WIDTH-1:0]     ns_arid,
  input  wire [NS_ADDR_WIDTH-1:0]   ns_araddr,
  output wire [NS_ID_WIDTH-1:0]     ns_rid,
  output wire [NS_DATA_WIDTH-1:0]   ns_rdata,
  input  wire [7:0] ns_awlen,
  input  wire [2:0] ns_awsize,
  input  wire [1:0] ns_awburst,
  input  wire       ns_awvalid,
  output wire       ns_awready,
  input  wire       ns_wlast,
  input  wire       ns_wvalid,
  output wire       ns_wready,
  output wire [1:0] ns_bresp,
  output wire       ns_bvalid,
  input  wire       ns_bready,
  input  wire [7:0] ns_arlen,
  input  wire [2:0] ns_arsize,
  input  wire [1:0] ns_arburst,
  input  wire       ns_arvalid,
  output wire       ns_arready,
  output wire [1:0] ns_rresp,
  output wire       ns_rlast,
  output wire       ns_rvalid,
  input  wire       ns_rready,

);

driver #(
  .HP_ADDR_WIDTH(HP_ADDR_WIDTH),
  .HP_DATA_WIDTH(HP_DATA_WIDTH),
  .LP_ADDR_WIDTH(LP_ADDR_WIDTH),
  .LP_DATA_WIDTH(LP_DATA_WIDTH),
  .NL_ADDR_WIDTH(NL_ADDR_WIDTH),
  .NL_DATA_WIDTH(NL_DATA_WIDTH),
  .NM_ADDR_WIDTH(NM_ADDR_WIDTH),
  .NM_DATA_WIDTH(NM_DATA_WIDTH),
  .NS_ID_WIDTH(NS_ID_WIDTH),
  .NS_ADDR_WIDTH(NS_ADDR_WIDTH),
  .NS_DATA_WIDTH(NS_DATA_WIDTH)
) driver_inst (
  .clk(clk),
  .rstn(rstn),
  .hp_awaddr  (hp_awaddr),
  .hp_wdata   (hp_wdata),
  .hp_wstrb   (hp_wstrb),
  .hp_araddr  (hp_araddr),
  .hp_rdata   (hp_rdata),
  .hp_awlen   (hp_awlen),
  .hp_awsize  (hp_awsize),
  .hp_awburst (hp_awburst),
  .hp_awvalid (hp_awvalid),
  .hp_awready (hp_awready),
  .hp_wlast   (hp_wlast),
  .hp_wvalid  (hp_wvalid),
  .hp_wready  (hp_wready),
  .hp_bresp   (hp_bresp),
  .hp_bvalid  (hp_bvalid),
  .hp_bready  (hp_bready),
  .hp_arlen   (hp_arlen),
  .hp_arsize  (hp_arsize),
  .hp_arburst (hp_arburst),
  .hp_arvalid (hp_arvalid),
  .hp_arready (hp_arready),
  .hp_rresp   (hp_rresp),
  .hp_rlast   (hp_rlast),
  .hp_rvalid  (hp_rvalid),
  .hp_rready  (hp_rready),
  .lp_awaddr  (lp_awaddr),
  .lp_wdata   (lp_wdata),
  .lp_wstrb   (lp_wstrb),
  .lp_araddr  (lp_araddr),
  .lp_rdata   (lp_rdata),
  .lp_awvalid (lp_awvalid),
  .lp_awready (lp_awready),
  .lp_wvalid  (lp_wvalid),
  .lp_wready  (lp_wready),
  .lp_bresp   (lp_bresp),
  .lp_bvalid  (lp_bvalid),
  .lp_bready  (lp_bready),
  .lp_arvalid (lp_arvalid),
  .lp_arready (lp_arready),
  .lp_rresp   (lp_rresp),
  .lp_rvalid  (lp_rvalid),
  .lp_rready  (lp_rready),
  .nl_awaddr  (nl_awaddr),
  .nl_wdata   (nl_wdata),
  .nl_wstrb   (nl_wstrb),
  .nl_araddr  (nl_araddr),
  .nl_rdata   (nl_rdata),
  .nl_awvalid (nl_awvalid),
  .nl_awready (nl_awready),
  .nl_wvalid  (nl_wvalid),
  .nl_wready  (nl_wready),
  .nl_bresp   (nl_bresp),
  .nl_bvalid  (nl_bvalid),
  .nl_bready  (nl_bready),
  .nl_arvalid (nl_arvalid),
  .nl_arready (nl_arready),
  .nl_rresp   (nl_rresp),
  .nl_rvalid  (nl_rvalid),
  .nl_rready  (nl_rready),
  .nm_awaddr  (nm_awaddr),
  .nm_wdata   (nm_wdata),
  .nm_wstrb   (nm_wstrb),
  .nm_araddr  (nm_araddr),
  .nm_rdata   (nm_rdata),
  .nm_awlen   (nm_awlen),
  .nm_awsize  (nm_awsize),
  .nm_awburst (nm_awburst),
  .nm_awvalid (nm_awvalid),
  .nm_awready (nm_awready),
  .nm_wlast   (nm_wlast),
  .nm_wvalid  (nm_wvalid),
  .nm_wready  (nm_wready),
  .nm_bresp   (nm_bresp),
  .nm_bvalid  (nm_bvalid),
  .nm_bready  (nm_bready),
  .nm_arlen   (nm_arlen),
  .nm_arsize  (nm_arsize),
  .nm_arburst (nm_arburst),
  .nm_arvalid (nm_arvalid),
  .nm_arready (nm_arready),
  .nm_rresp   (nm_rresp),
  .nm_rlast   (nm_rlast),
  .nm_rvalid  (nm_rvalid),
  .nm_rready  (nm_rready),
  .ns_awid    (ns_awid),
  .ns_awaddr  (ns_awaddr),
  .ns_wdata   (ns_wdata),
  .ns_wstrb   (ns_wstrb),
  .ns_bid     (ns_bid),
  .ns_arid    (ns_arid),
  .ns_araddr  (ns_araddr),
  .ns_rid     (ns_rid),
  .ns_rdata   (ns_rdata),
  .ns_awlen   (ns_awlen),
  .ns_awsize  (ns_awsize),
  .ns_awburst (ns_awburst),
  .ns_awvalid (ns_awvalid),
  .ns_awready (ns_awready),
  .ns_wlast   (ns_wlast),
  .ns_wvalid  (ns_wvalid),
  .ns_wready  (ns_wready),
  .ns_bresp   (ns_bresp),
  .ns_bvalid  (ns_bvalid),
  .ns_bready  (ns_bready),
  .ns_arlen   (ns_arlen),
  .ns_arsize  (ns_arsize),
  .ns_arburst (ns_arburst),
  .ns_arvalid (ns_arvalid),
  .ns_arready (ns_arready),
  .ns_rresp   (ns_rresp),
  .ns_rlast   (ns_rlast),
  .ns_rvalid  (ns_rvalid),
  .ns_rready  (ns_rready),

);

endmodule