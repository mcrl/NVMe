`timescale 1ps / 1ps

module top (
  // System Interface
  input sys_clk_p,
  input sys_clk_n,
  input sys_rst_n,

  // PCIe serial 
  output pci_exp_txp,
  output pci_exp_txn,
  input pci_exp_rxp,
  input pci_exp_rxn
);


endmodule
